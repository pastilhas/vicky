module qoi

fn encode() {
}
